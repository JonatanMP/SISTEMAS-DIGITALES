module andcompuerta ( input a, b, 
output v);

assign v=(a&b);

endmodule   