module tratamiento de datos ( 
    input reg datokey,
    output reg cont

    
);
 reg dato1, dato;
 count = 0;

 always @(posedge clkot) begin
    count = 
    if (dato1 == 4'b0000 && dato <= 4'b0000 ) begin
        count = count + 1;
    end
    else count = count
        
 end

//  always @(posedge clkot) begin //contaor con la salida del clock dividido para control de displays 
//     ct <= ct+2'd1;    
//     if (ct == 2'b11)
//     ct <= 2'b00;
//     else
//     ct <= ct + 1;
  
// end


always @(posedge tecla del teclado precionada and  contador de primer datos) begin


    
end

endmodule //tratamiento de datos